// fp32_div.v
//
// Verilog RTL for a 32-bit (single-precision) floating-point divider.
//
// Operation: result = a / b
//
// Format (IEEE 754 single-precision):
// [31]   : Sign bit
// [30:23]: 8-bit exponent (bias of 127)
// [22:0] : 23-bit mantissa
//
// Features:
// - Fixed-latency 26-stage pipelined architecture.
// - Uses a pipelined restoring division algorithm for the mantissa.
// - Handles normalized and denormalized numbers.
// - Handles special cases: NaN, Infinity, Zero, and Division by Zero.
// - Truncates the result.

module fp32_div (
    input clk,
    input rst_n,
    input  [31:0] a,
    input  [31:0] b,
    output [31:0] result
);

    // Latency of the divider core = 24 cycles (23 mantissa bits + 1 integer bit)
    localparam DIV_LATENCY = 24;
    localparam TOTAL_LATENCY = DIV_LATENCY + 1;

    //----------------------------------------------------------------
    // Stage 1: Unpack and Handle Special Cases
    //----------------------------------------------------------------
    
    wire        sign_a = a[31];
    wire [ 7:0] exp_a  = a[30:23];
    wire [22:0] mant_a = a[22:0];

    wire        sign_b = b[31];
    wire [ 7:0] exp_b  = b[30:23];
    wire [22:0] mant_b = b[22:0];

    // Detect special values
    wire is_nan_a = (exp_a == 8'hFF) && (mant_a != 0);
    wire is_inf_a = (exp_a == 8'hFF) && (mant_a == 0);
    wire is_zero_a = (exp_a == 0) && (mant_a == 0);

    wire is_nan_b = (exp_b == 8'hFF) && (mant_b != 0);
    wire is_inf_b = (exp_b == 8'hFF) && (mant_b == 0);
    wire is_zero_b = (exp_b == 0) && (mant_b == 0);

    // Add implicit leading bit
    wire [23:0] full_mant_a = {(exp_a != 0), mant_a};
    wire [23:0] full_mant_b = {(exp_b != 0), mant_b};

    wire [ 8:0] eff_exp_a = (exp_a == 0) ? 1 : exp_a;
    wire [ 8:0] eff_exp_b = (exp_b == 0) ? 1 : exp_b;

    // Stage 1 Pipeline Registers
    reg         s1_special_case;
    reg  [31:0] s1_special_result;
    reg  signed [8:0] s1_exp_res;
    reg         s1_sign_res;
    reg  [46:0] s1_dividend; // For (mant_a << 23)
    reg  [23:0] s1_divisor;

    always @(posedge clk) begin
        if (!rst_n) begin
            s1_special_case <= 1'b0;
            s1_special_result <= 32'b0;
            s1_exp_res <= 9'b0;
            s1_sign_res <= 1'b0;
            s1_dividend <= 47'b0;
            s1_divisor <= 24'b0;
        end else begin
            // Default path for normal operation
            s1_special_case <= 1'b0;
            s1_dividend <= {full_mant_a, 23'b0};
            s1_divisor <= full_mant_b;
            s1_sign_res <= sign_a ^ sign_b;

            s1_exp_res <= eff_exp_a - eff_exp_b + 127;

            // Handle special cases
            if (is_nan_a || is_nan_b || (is_inf_a && is_inf_b) || (is_zero_a && is_zero_b)) begin
                s1_special_case <= 1'b1;
                s1_special_result <= 32'h7FC00001; // qNaN
            end else if (is_inf_a || is_zero_b) begin
                s1_special_case <= 1'b1;
                s1_special_result <= {sign_a ^ sign_b, 8'hFF, 23'b0}; // Infinity
            end else if (is_zero_a || is_inf_b) begin
                s1_special_case <= 1'b1;
                s1_special_result <= {sign_a ^ sign_b, 31'b0}; // Zero
            end
        end
    end

    //----------------------------------------------------------------
    // Pipelined Divider Core (24 Stages)
    //----------------------------------------------------------------
    
    // Arrays of registers to pipeline the division state
    reg  [24:0] rem_pipe      [0:DIV_LATENCY];
    reg  [46:0] dividend_pipe [0:DIV_LATENCY];
    reg  [23:0] divisor_pipe  [0:DIV_LATENCY];
    reg  [23:0] quotient_pipe [0:DIV_LATENCY];

    // Initialize first stage of the divider pipeline
    always @(posedge clk) begin
        if (!rst_n) begin
            rem_pipe[0] <= 25'b0;
            dividend_pipe[0] <= 47'b0;
            divisor_pipe[0] <= 24'b0;
            quotient_pipe[0] <= 24'b0;
        end else begin
            rem_pipe[0] <= 25'b0;
            dividend_pipe[0] <= s1_dividend;
            divisor_pipe[0] <= s1_divisor;
            quotient_pipe[0] <= 24'b0;
        end
    end

    // Generate the divider stages
    genvar i;
    generate
        for (i = 0; i < DIV_LATENCY; i = i + 1) begin : div_stages
            // Combinational logic for one stage of restoring division
            wire [24:0] shifted_rem = {rem_pipe[i][23:0], dividend_pipe[i][46]};
            wire [24:0] sub_res = shifted_rem - {1'b0, divisor_pipe[i]};
            wire q_bit = ~sub_res[24];

            // Register the results for the next stage
            always @(posedge clk) begin
                if(!rst_n) begin
                    rem_pipe[i+1] <= 25'b0;
                    dividend_pipe[i+1] <= 47'b0;
                    divisor_pipe[i+1] <= 24'b0;
                    quotient_pipe[i+1] <= 24'b0;
                end else begin
                    rem_pipe[i+1] <= q_bit ? sub_res : shifted_rem;
                    dividend_pipe[i+1] <= dividend_pipe[i] << 1;
                    divisor_pipe[i+1] <= divisor_pipe[i];
                    quotient_pipe[i+1] <= {quotient_pipe[i][22:0], q_bit};
                end
            end
        end
    endgenerate

    // Pipeline to carry special flags and results alongside the divider
    reg [TOTAL_LATENCY:0] special_case_pipe;
    reg [31:0] special_result_pipe [TOTAL_LATENCY:0];
    reg signed [8:0] exp_res_pipe [TOTAL_LATENCY:0];
    reg sign_res_pipe [TOTAL_LATENCY:0];

    always @(posedge clk) begin
        if(!rst_n) begin
            special_case_pipe[0] <= 1'b0;
            special_result_pipe[0] <= 32'b0;
            exp_res_pipe[0] <= 9'b0;
            sign_res_pipe[0] <= 1'b0;
        end else begin
            special_case_pipe[0] <= s1_special_case;
            special_result_pipe[0] <= s1_special_result;
            exp_res_pipe[0] <= s1_exp_res;
            sign_res_pipe[0] <= s1_sign_res;
        end
    end
    
    generate
        for(i=0; i<TOTAL_LATENCY; i=i+1) begin : prop_pipe
            always @(posedge clk) begin
                if(!rst_n) begin
                    special_case_pipe[i+1] <= 1'b0;
                    special_result_pipe[i+1] <= 32'b0;
                    exp_res_pipe[i+1] <= 9'b0;
                    sign_res_pipe[i+1] <= 1'b0;
                end else begin
                    special_case_pipe[i+1] <= special_case_pipe[i];
                    special_result_pipe[i+1] <= special_result_pipe[i];
                    exp_res_pipe[i+1] <= exp_res_pipe[i];
                    sign_res_pipe[i+1] <= sign_res_pipe[i];
                end
            end
        end
    endgenerate

    //----------------------------------------------------------------
    // Final Stage: Normalize and Pack
    //----------------------------------------------------------------
    
    // Result of the mantissa division
    wire [23:0] final_quotient = quotient_pipe[DIV_LATENCY];
    
    // Normalize the mantissa and adjust exponent
    reg  signed [ 8:0] final_exp;
    reg         [22:0] final_mant;
    
    always @(*) begin
        // The division of two normalized mantissas (1.f / 1.f) gives a result
        // in the range [0.5, 2.0).
        // If the result is < 1.0 (quotient[23]==0), we must normalize left.
        if(!final_quotient[23]) begin
            final_exp = exp_res_pipe[TOTAL_LATENCY] - 1;
            final_mant = final_quotient[22:0] << 1; 
        end else begin
            final_exp = exp_res_pipe[TOTAL_LATENCY];
            final_mant = final_quotient[22:0];
        end
    end
    
    // Handle final exponent overflow/underflow
    reg  [ 7:0] out_exp;
    reg  [22:0] out_mant;
    
    always @(*) begin
        out_exp = final_exp[7:0];
        out_mant = final_mant;
        
        if (final_exp >= 255) begin // Overflow -> Inf
            out_exp = 8'hFF;
            out_mant = 23'b0;
        end else if (final_exp <= 0) begin // Underflow -> Denormalized or Zero
            out_mant = ({1'b1, final_mant}) >> (1 - final_exp);
            out_exp = 8'b0;
        end
    end
    
    // Final registered output
    reg  [31:0] result_reg;
    always @(posedge clk) begin
        if (!rst_n) begin
            result_reg <= 32'b0;
        end else begin
            if (special_case_pipe[TOTAL_LATENCY]) begin
                result_reg <= special_result_pipe[TOTAL_LATENCY];
            end else if (out_exp == 0 && out_mant == 0) begin
                result_reg <= {sign_res_pipe[TOTAL_LATENCY], 31'b0};
            end else begin
                result_reg <= {sign_res_pipe[TOTAL_LATENCY], out_exp, out_mant};
            end
        end
    end
    
    assign result = result_reg;

endmodule
